module subArray #(

//-------------------Shared Parameters with controller  
   parameter OPERATION_WIDTH=1,  //for ALU with two operations
   parameter SRC_WIDTH=2, 
   parameter NUM_OF_COL_IN_ROW=64,
   parameter NUM_ROW_IN_SUBARRAY=1024,
   parameter ROW_CYCLE=50, //ns
   parameter SHIFT_CYCLE=6, //ns 
   parameter NUMBER_OF_WAIT_CYCLE_FOR_ROW_LOAD=9,  //$ceil(ROW_CYCLE/SHIFT_CYCLE),
   parameter WAIT_CYCLE_WIDTH=4   ,        //$ceil($clog2(NUMBER_OF_WAIT_CYCLE_FOR_ROW_LOAD)),
   parameter COL_COUNTER_WIDTH=6,      //$ceil($clog2(NUM_OF_COL_IN_ROW)),
   parameter ROW_ADR_WIDTH=10,// $ceil($clog2(NUM_ROW_IN_SUBARRAY)),
   parameter COMMAND_WIDTH=4,
   parameter GOLOBAL_DATA_BUS_WIDTH=32,
   parameter OUT_SRC_WIDTH=1,
//------OPCODE ENCODING
  parameter ADD_OPCODE=0,
  parameter MULT_OPCODE=1,
//-----------SRC SELCTION ENCODING
   parameter SRC_ROW1=0,
   parameter SRC_ROW2=1,
   parameter SRC_GLLOBAL_BUS=2,
   parameter SRC_TEMP_REG_A=3,
   parameter SRC_TEMP_REG_B=4,
   parameter SRC_TEMP_REG_C=5,
   parameter SRC_TEMP_ADDER_OUT=6,
   parameter SRC_TEMP_MULTIPLIER_OUT=7,
//---------------READ_WRITE_ENCODING
   parameter READ=0,
   parameter WRITE=1,
   //-------------Extra parameters to be removed ----------------------
   parameter addedToKeepCommaLess=0

)(
   //-------------Input Ports-----------------------------
   input logic clk,           // clock
   input logic reset,         // Active high, syn reset
   input logic start,
   input logic valid_command, // Request 0
   input logic [ ROW_ADR_WIDTH-1:0] row_addr,
   input logic [ COMMAND_WIDTH-1:0] command,
   input logic [GOLOBAL_DATA_BUS_WIDTH-1:0] global_data_bus,
   input logic [NUM_OF_COL_IN_ROW-1:0] [GOLOBAL_DATA_BUS_WIDTH-1:0] rowFromSubarray,
   //output ports
   output logic [NUM_OF_COL_IN_ROW-1:0] [GOLOBAL_DATA_BUS_WIDTH-1:0] rowToSubarray
   );

//---------------------Internal Variables
   //Controller's ports
   logic [0:0] shift1;
   logic [0:0] shift2;
   logic [0:0] shift3;
   logic [0:0] shiftDir1_read_or_write;
   logic [0:0] shiftDir2_read_or_write;
   logic [0:0] shiftDir3_read_or_write;
   logic [OPERATION_WIDTH-1:0] opCode1;
   logic [OPERATION_WIDTH-1:0] opCode2;
   logic [SRC_WIDTH-1:0] src1Op1;
   logic [SRC_WIDTH-1:0] src2Op1;
   logic [SRC_WIDTH-1:0] src1Op2;
   logic [SRC_WIDTH-1:0] src2Op2;
   logic read_or_write;
   logic row1_active;
   logic row2_active;
   logic row3_active;

   logic load_temp_regA;
   logic load_temp_regB;
   logic load_temp_regC;
   
//Shift Registers signal
   logic [NUM_OF_COL_IN_ROW-1:0] [GOLOBAL_DATA_BUS_WIDTH-1:0] outputRow1;
   logic [NUM_OF_COL_IN_ROW-1:0] [GOLOBAL_DATA_BUS_WIDTH-1:0] outputRow2;
   logic [NUM_OF_COL_IN_ROW-1:0] [GOLOBAL_DATA_BUS_WIDTH-1:0] outputRow3;
//------------------temp registers
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0]  temp_regA;
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0]  temp_regB;
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0]  temp_regC;

//---------------Adder  input signals
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0] adder_input1;
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0] adder_input2 ;
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0] adder_output1;
   logic [SRC_WIDTH-1:0] src1Adder;
   logic [SRC_WIDTH-1:0] src2Adder;
   logic [SRC_WIDTH-1:0] src1Multiplier;
   logic [SRC_WIDTH-1:0] src2Multiplier;
//---------------Signals automatically generated by mpdole instanciation   
   //logic equalFlag;
   //logic lessFlag;

//--------------multiplier input signals
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0] multiplier_input1;
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0] multiplier_input2 ;
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0] multiplier_output1;
//--------------------------------------Row signals
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0] inputColumnRow1;
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0] inputColumnRow2 ;
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0] inputColumnRow3;

   logic [GOLOBAL_DATA_BUS_WIDTH-1:0]  outputColumnRow1;
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0] outputColumnRow2 ;
   logic [GOLOBAL_DATA_BUS_WIDTH-1:0] outputColumnRow3;

   logic loadRow1;
   logic loadRow2;
   logic loadRow3;

//------------------------------------

multiplier#(
.GOLOBAL_DATA_BUS_WIDTH(GOLOBAL_DATA_BUS_WIDTH))
 multiplier_instance1(
.input1(multiplier_input1),
.input2(multiplier_input2),
.output1(multiplier_output1)
);
//assign rowToSubarray[1]=multiplier_output1; //debug line 

//--------------------------------------
adder#(
.GOLOBAL_DATA_BUS_WIDTH(GOLOBAL_DATA_BUS_WIDTH)) 
 adder_instance1(
.input1(adder_input1),
.input2(adder_input2),
.output1(adder_output1),
.equalFlag(equalFlag),
.lessFlag(lessFlag)
);
//assign rowToSubarray[2]=multiplier_output1; //debug line
//-----------------------------------------------------
controller_programmable#(
  .OPERATION_WIDTH(OPERATION_WIDTH),  //for ALU with two operations
  .SRC_WIDTH(SRC_WIDTH), 
   .NUM_OF_COL_IN_ROW(NUM_OF_COL_IN_ROW),
   .NUM_ROW_IN_SUBARRAY(NUM_ROW_IN_SUBARRAY),
   .NUMBER_OF_WAIT_CYCLE_FOR_ROW_LOAD(NUMBER_OF_WAIT_CYCLE_FOR_ROW_LOAD),
   .WAIT_CYCLE_WIDTH(WAIT_CYCLE_WIDTH),
   .COL_COUNTER_WIDTH(COL_COUNTER_WIDTH),
   .ROW_ADR_WIDTH(ROW_ADR_WIDTH),
   .COMMAND_WIDTH(COMMAND_WIDTH),
   .GOLOBAL_DATA_BUS_WIDTH(GOLOBAL_DATA_BUS_WIDTH),
   .OUT_SRC_WIDTH(OUT_SRC_WIDTH)

)
 controller_instance1
(
   .clk(clk), 
   .reset(reset), .start(start),.valid_command(valid_command),   
   .row_addr(row_addr),
   .command(command),
   .global_data_bus(global_data_bus), //TODO: implement systolic GDls here
  .adder_equal_flag(equalFlag),
   .adder_less_flag(lessFlag),
   //-----------------
//---------------------
   .shift1(shift1),
   .shift2(shift2),
   .shift3(shift3),
   .shiftDir1_read_or_write(shiftDir1_read_or_write),
   .shiftDir2_read_or_write(shiftDir2_read_or_write),
   .shiftDir3_read_or_write(shiftDir3_read_or_write),
   .opCode1(opCode1),
   .opCode2(opCode2),
   .src1Op1(src1Op1),
   .src2Op1(src2Op1),
   .src1Op2(src1Op2),
   .src2Op2(src2Op2),
   .read_or_write(read_or_write),
   .row1_active(row1_active),
   .row2_active(row2_active),
   .row3_active(row3_active),
   .load_temp_regA(load_temp_regA),
   .load_temp_regB(load_temp_regB),
   .load_temp_regC(load_temp_regC),
   .pc(pc),
   .outShiftValueSrc(outShiftValueSrc)
   );


//-----------------------------------
row_wide_shifter #(
.GOLOBAL_DATA_BUS_WIDTH(GOLOBAL_DATA_BUS_WIDTH),
.NUM_OF_COL_IN_ROW(NUM_OF_COL_IN_ROW)
)row_wide_shifter_instance1
(
.clk(clk),
.loadRow(loadRow1),
.inputRow(rowFromSubarray),
.inputColumn(inputColumnRow1),
.shiftSignal(shift1),
.shiftDir_read_or_write(shiftDir1_read_or_write), //1 right, 0 
//-------
.outputRow(outputRow1),
.outputColumn(outputColumnRow1)
);
//---------------------------------
row_wide_shifter #(
.GOLOBAL_DATA_BUS_WIDTH(GOLOBAL_DATA_BUS_WIDTH),
.NUM_OF_COL_IN_ROW(NUM_OF_COL_IN_ROW)
)row_wide_shifter_instance2
(
.clk(clk),
.loadRow(loadRow2),
.inputRow(rowFromSubarray),
.inputColumn(inputColumnRow2),
.shiftSignal(shift2),
.shiftDir_read_or_write(shiftDir2_read_or_write), //read 0, write 1
//-------
.outputRow(outputRow2),
.outputColumn(outputColumnRow2)
);
//----------------------------------
row_wide_shifter #(
.GOLOBAL_DATA_BUS_WIDTH(GOLOBAL_DATA_BUS_WIDTH),
.NUM_OF_COL_IN_ROW(NUM_OF_COL_IN_ROW)
)row_wide_shifter_instance3
(
.clk(clk),
.loadRow(loadRow3),
.inputRow(rowFromSubarray),
.inputColumn(inputColumnRow3),
.shiftSignal(shift3),
.shiftDir_read_or_write(shiftDir3_read_or_write), //read 0, write 1
//-------
.outputRow(outputRow3),
.outputColumn(outputColumnRow3)
);
//--------------------------------------Assigning input and output of signals
  assign inputColumnRow1 = outShiftValueSrc ? adder_output1:  multiplier_output1;
  assign inputColumnRow2 = outShiftValueSrc ? adder_output1:  multiplier_output1;
  assign inputColumnRow3 = outShiftValueSrc ? adder_output1:  multiplier_output1;
//-------------------------------------
   assign loadRow1 = row1_active & (read_or_write==READ);
   assign loadRow2 = row2_active & (read_or_write==READ);
   assign loadRow3 = row3_active & (read_or_write==READ);
//-------------------------------------
   assign src1Adder= (opCode1 == ADD_OPCODE) ? src1Op1 : src1Op2; //TODO: assume that ALU has only two operations
   assign src2Adder= (opCode1 == ADD_OPCODE) ? src2Op1 : src2Op2;
   assign src1Multiplier =(opCode1 == MULT_OPCODE) ? src1Op1 : src1Op2;
   assign src2Multiplier =(opCode1 == MULT_OPCODE) ? src2Op1 : src2Op2;
//------------------------------------
assign rowToSubarray=read_or_write ?(row1_active ? (outputRow1):(row2_active ?outputRow2:outputRow3 )):(0); //debug commented
/*
always @(*) begin
  
  case({{read_or_write},{row1_active},{row1_active},{row1_active}})
     4'b1100:begin
   	rowToSubarray<=outputRow1;
     end
     4'b1010:begin
   	rowToSubarray<=outputRow2;
     end
     4'b1001:begin
   	 rowToSubarray<=outputRow3;
     end
     default:begin
         rowToSubarray<=0;
     end
    endcase;
  
end
*/
//------------------------
always_comb begin
  
  case(src1Adder) 
    SRC_ROW1: begin
   		adder_input1<=outputColumnRow1;
    end	
    SRC_ROW2: begin
		adder_input1<=outputColumnRow2;
    end
    SRC_GLLOBAL_BUS: begin
		adder_input1<=global_data_bus;
    end
    SRC_TEMP_REG_A: begin
		adder_input1<=temp_regA;
    end
    SRC_TEMP_REG_B: begin
		adder_input1<=temp_regB;
    end
    SRC_TEMP_REG_C: begin
	       adder_input1<=temp_regC;
    end
    SRC_TEMP_ADDER_OUT: begin
		adder_input1<=adder_output1;
     end
    SRC_TEMP_MULTIPLIER_OUT: begin
		adder_input1<=multiplier_output1;
     end
     default:begin
                 adder_input1<=0;
    end
    endcase;
  
end

always_comb begin
  
  case(src2Adder) 
    SRC_ROW1: begin
   		adder_input2<=outputColumnRow1;
    end	
    SRC_ROW2: begin
		adder_input2<=outputColumnRow2;
    end
    SRC_GLLOBAL_BUS: begin
		adder_input2<=global_data_bus;
    end
    SRC_TEMP_REG_A: begin
		adder_input2<=temp_regA;
    end
    SRC_TEMP_REG_B: begin
		adder_input2<=temp_regB;
    end
    SRC_TEMP_REG_C: begin
	       adder_input2<=temp_regC;
    end
    SRC_TEMP_ADDER_OUT: begin
		adder_input2<=adder_output1;
     end
    SRC_TEMP_MULTIPLIER_OUT: begin
		adder_input2<=multiplier_output1;
     end
     default:begin
                 adder_input2<=0;
    end
    endcase;
 
  
end
//--------------------

always_comb begin
  
  case(src1Multiplier) 
    SRC_ROW1: begin
   		multiplier_input1<=outputColumnRow1;
    end	
    SRC_ROW2: begin
		multiplier_input1<=outputColumnRow2;
    end
    SRC_GLLOBAL_BUS: begin
		multiplier_input1<=global_data_bus;
    end
    SRC_TEMP_REG_A: begin
		multiplier_input1<=temp_regA;
    end
    SRC_TEMP_REG_B: begin
		multiplier_input1<=temp_regB;
    end
    SRC_TEMP_REG_C: begin
	       multiplier_input1<=temp_regC;
    end
    SRC_TEMP_ADDER_OUT: begin
		multiplier_input1<=adder_output1;
     end
    SRC_TEMP_MULTIPLIER_OUT: begin
		multiplier_input1<=multiplier_output1;
     end
     default:begin
                 multiplier_input1<=0;
    end
    endcase;
 
  
end
always_comb begin
  
  case(src2Multiplier) 
    SRC_ROW1: begin
   		multiplier_input2<=outputColumnRow1;
    end	
    SRC_ROW2: begin
		multiplier_input2<=outputColumnRow2;
    end
    SRC_GLLOBAL_BUS: begin
		multiplier_input2<=outputColumnRow3;
    end
    SRC_TEMP_REG_A: begin
		multiplier_input2<=temp_regA;
    end
    SRC_TEMP_REG_B: begin
		multiplier_input2<=temp_regB;
    end
    SRC_TEMP_REG_C: begin
	       multiplier_input2<=temp_regC;
    end
    SRC_TEMP_ADDER_OUT: begin
		multiplier_input2<=adder_output1;
     end
    SRC_TEMP_MULTIPLIER_OUT: begin
		multiplier_input2<=multiplier_output1;
     end
     default:begin
                 multiplier_input2<=0;
    end
    endcase;
 
  
end


always @ (posedge clk or posedge reset ) begin : TEMP_REG_A_MAINTAIN
	if (reset) begin
		temp_regA<=0;
	end else begin
		if (load_temp_regA) begin
			temp_regA<=global_data_bus;
		end
	end 
end
always @ (posedge clk or posedge reset) begin : TEMP_REG_B_MAINTAIN
	if (reset) begin
		temp_regB<=0;
	end else begin
		if (load_temp_regB) begin
			temp_regB<=global_data_bus;
		end
	end 
end
always @ (posedge clk or posedge reset ) begin : TEMP_REG_C_MAINTAIN
	if (reset) begin
		temp_regC<=0;
	end else begin
		if (load_temp_regC) begin
			temp_regC<=global_data_bus;
		end
	end 
end

endmodule // End of Module controller




